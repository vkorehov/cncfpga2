`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:12:59 05/22/2014 
// Design Name: 
// Module Name:    cnc_top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cnc_top(
    inout [31:0] AD,
    inout [3:0] CBE_N,
	 inout PAR,
    inout FRAME_N,
    inout TRDY_N,
    inout IRDY_N,
    inout STOP_N,
    inout DEVSEL_N,
    input IDSEL,
    output INTA_N,
    inout PERR_N,
    inout SERR_N,
    output REQ_N,
    input GNT_N,
    input RST_N,
    input PCLK,
    output PING_DONE,
    input PING_REQ
    );

// I/O structure instantiations

IOBUF_PCI33_5 XPCI_ADB31 (.O(AD_I31),.IO(AD[31]),.I(AD_OUT31),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB30 (.O(AD_I30),.IO(AD[30]),.I(AD_OUT30),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB29 (.O(AD_I29),.IO(AD[29]),.I(AD_OUT29),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB28 (.O(AD_I28),.IO(AD[28]),.I(AD_OUT28),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB27 (.O(AD_I27),.IO(AD[27]),.I(AD_OUT27),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB26 (.O(AD_I26),.IO(AD[26]),.I(AD_OUT26),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB25 (.O(AD_I25),.IO(AD[25]),.I(AD_OUT25),.T(OE_AD3_N   ));
IOBUF_PCI33_5 XPCI_ADB24 (.O(AD_I24),.IO(AD[24]),.I(AD_OUT24),.T(OE_AD3_N   ));

IOBUF_PCI33_5 XPCI_ADB23 (.O(AD_I23),.IO(AD[23]),.I(AD_OUT23),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB22 (.O(AD_I22),.IO(AD[22]),.I(AD_OUT22),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB21 (.O(AD_I21),.IO(AD[21]),.I(AD_OUT21),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB20 (.O(AD_I20),.IO(AD[20]),.I(AD_OUT20),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB19 (.O(AD_I19),.IO(AD[19]),.I(AD_OUT19),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB18 (.O(AD_I18),.IO(AD[18]),.I(AD_OUT18),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB17 (.O(AD_I17),.IO(AD[17]),.I(AD_OUT17),.T(OE_AD2_N  ));
IOBUF_PCI33_5 XPCI_ADB16 (.O(AD_I16),.IO(AD[16]),.I(AD_OUT16),.T(OE_AD2_N  ));

IOBUF_PCI33_5 XPCI_ADB15 (.O(AD_I15),.IO(AD[15]),.I(AD_OUT15),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB14 (.O(AD_I14),.IO(AD[14]),.I(AD_OUT14),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB13 (.O(AD_I13),.IO(AD[13]),.I(AD_OUT13),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB12 (.O(AD_I12),.IO(AD[12]),.I(AD_OUT12),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB11 (.O(AD_I11),.IO(AD[11]),.I(AD_OUT11),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB10 (.O(AD_I10),.IO(AD[10]),.I(AD_OUT10),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB9  (.O(AD_I9 ),.IO(AD[9 ]),.I(AD_OUT9 ),.T(OE_AD1_N  ));
IOBUF_PCI33_5 XPCI_ADB8  (.O(AD_I8 ),.IO(AD[8 ]),.I(AD_OUT8 ),.T(OE_AD1_N  ));

IOBUF_PCI33_5 XPCI_ADB7  (.O(AD_I7 ),.IO(AD[7 ]),.I(AD_OUT7 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB6  (.O(AD_I6 ),.IO(AD[6 ]),.I(AD_OUT6 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB5  (.O(AD_I5 ),.IO(AD[5 ]),.I(AD_OUT5 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB4  (.O(AD_I4 ),.IO(AD[4 ]),.I(AD_OUT4 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB3  (.O(AD_I3 ),.IO(AD[3 ]),.I(AD_OUT3 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB2  (.O(AD_I2 ),.IO(AD[2 ]),.I(AD_OUT2 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB1  (.O(AD_I1 ),.IO(AD[1 ]),.I(AD_OUT1 ),.T(OE_AD0_N   ));
IOBUF_PCI33_5 XPCI_ADB0  (.O(AD_I0 ),.IO(AD[0 ]),.I(AD_OUT0 ),.T(OE_AD0_N   ));
// input flipflops
FDPE XPCI_ADIQ31 (.Q(AD31),.D(AD_I31),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ30 (.Q(AD30),.D(AD_I30),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ29 (.Q(AD29),.D(AD_I29),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ28 (.Q(AD28),.D(AD_I28),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ27 (.Q(AD27),.D(AD_I27),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ26 (.Q(AD26),.D(AD_I26),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ25 (.Q(AD25),.D(AD_I25),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ24 (.Q(AD24),.D(AD_I24),.C(CLK),.CE(1'b1),.PRE(RST));

FDPE XPCI_ADIQ23 (.Q(AD23),.D(AD_I23),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ22 (.Q(AD22),.D(AD_I22),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ21 (.Q(AD21),.D(AD_I21),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ20 (.Q(AD20),.D(AD_I20),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ19 (.Q(AD19),.D(AD_I19),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ18 (.Q(AD18),.D(AD_I18),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ17 (.Q(AD17),.D(AD_I17),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ16 (.Q(AD16),.D(AD_I16),.C(CLK),.CE(1'b1),.PRE(RST));

FDPE XPCI_ADIQ15 (.Q(AD15),.D(AD_I15),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ14 (.Q(AD14),.D(AD_I14),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ13 (.Q(AD13),.D(AD_I13),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ12 (.Q(AD12),.D(AD_I12),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ11 (.Q(AD11),.D(AD_I11),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ10 (.Q(AD10),.D(AD_I10),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ9  (.Q(AD9 ),.D(AD_I9 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ8  (.Q(AD8 ),.D(AD_I8 ),.C(CLK),.CE(1'b1),.PRE(RST));

FDPE XPCI_ADIQ7  (.Q(AD7 ),.D(AD_I7 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ6  (.Q(AD6 ),.D(AD_I6 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ5  (.Q(AD5 ),.D(AD_I5 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ4  (.Q(AD4 ),.D(AD_I4 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ3  (.Q(AD3 ),.D(AD_I3 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ2  (.Q(AD2 ),.D(AD_I2 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ1  (.Q(AD1 ),.D(AD_I1 ),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_ADIQ0  (.Q(AD0 ),.D(AD_I0 ),.C(CLK),.CE(1'b1),.PRE(RST));
// output flipflops
FDE XPCI_ADOQ31 (.Q(AD_OUT31),.D(AD_O31),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ30 (.Q(AD_OUT30),.D(AD_O30),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ29 (.Q(AD_OUT29),.D(AD_O29),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ28 (.Q(AD_OUT28),.D(AD_O28),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ27 (.Q(AD_OUT27),.D(AD_O27),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ26 (.Q(AD_OUT26),.D(AD_O26),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ25 (.Q(AD_OUT25),.D(AD_O25),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ24 (.Q(AD_OUT24),.D(AD_O24),.C(CLK),.CE(PCI_CE));

FDE XPCI_ADOQ23 (.Q(AD_OUT23),.D(AD_O23),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ22 (.Q(AD_OUT22),.D(AD_O22),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ21 (.Q(AD_OUT21),.D(AD_O21),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ20 (.Q(AD_OUT20),.D(AD_O20),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ19 (.Q(AD_OUT19),.D(AD_O19),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ18 (.Q(AD_OUT18),.D(AD_O18),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ17 (.Q(AD_OUT17),.D(AD_O17),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ16 (.Q(AD_OUT16),.D(AD_O16),.C(CLK),.CE(PCI_CE));

FDE XPCI_ADOQ15 (.Q(AD_OUT15),.D(AD_O15),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ14 (.Q(AD_OUT14),.D(AD_O14),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ13 (.Q(AD_OUT13),.D(AD_O13),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ12 (.Q(AD_OUT12),.D(AD_O12),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ11 (.Q(AD_OUT11),.D(AD_O11),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ10 (.Q(AD_OUT10),.D(AD_O10),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ9  (.Q(AD_OUT9 ),.D(AD_O9 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ8  (.Q(AD_OUT8 ),.D(AD_O8 ),.C(CLK),.CE(PCI_CE));

FDE XPCI_ADOQ7  (.Q(AD_OUT7 ),.D(AD_O7 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ6  (.Q(AD_OUT6 ),.D(AD_O6 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ5  (.Q(AD_OUT5 ),.D(AD_O5 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ4  (.Q(AD_OUT4 ),.D(AD_O4 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ3  (.Q(AD_OUT3 ),.D(AD_O3 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ2  (.Q(AD_OUT2 ),.D(AD_O2 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ1  (.Q(AD_OUT1 ),.D(AD_O1 ),.C(CLK),.CE(PCI_CE));
FDE XPCI_ADOQ0  (.Q(AD_OUT0 ),.D(AD_O0 ),.C(CLK),.CE(PCI_CE));

IOBUF_PCI33_5 XPCI_CBB3 (.O(CBE_I3),.IO(CBE_N[3]),.I(CBE_OUT3),.T(OE_CBE_N  ));
IOBUF_PCI33_5 XPCI_CBB2 (.O(CBE_I2),.IO(CBE_N[2]),.I(CBE_OUT2),.T(OE_CBE_N  ));
IOBUF_PCI33_5 XPCI_CBB1 (.O(CBE_I1),.IO(CBE_N[1]),.I(CBE_OUT1),.T(OE_CBE_N  ));
IOBUF_PCI33_5 XPCI_CBB0 (.O(CBE_I0),.IO(CBE_N[0]),.I(CBE_OUT0),.T(OE_CBE_N  ));
// input flipflops
FDPE XPCI_CBIQ3 (.Q(CBE3),.D(CBE_I3),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_CBIQ2 (.Q(CBE2),.D(CBE_I2),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_CBIQ1 (.Q(CBE1),.D(CBE_I1),.C(CLK),.CE(1'b1),.PRE(RST));
FDPE XPCI_CBIQ0 (.Q(CBE0),.D(CBE_I0),.C(CLK),.CE(1'b1),.PRE(RST));
// output flipflops
FDE XPCI_CBOQ3 (.Q(CBE_OUT3),.D(CBE_O3),.C(CLK),.CE(PCI_CE));
FDE XPCI_CBOQ2 (.Q(CBE_OUT2),.D(CBE_O2),.C(CLK),.CE(PCI_CE));
FDE XPCI_CBOQ1 (.Q(CBE_OUT1),.D(CBE_O1),.C(CLK),.CE(PCI_CE));
FDE XPCI_CBOQ0 (.Q(CBE_OUT0),.D(CBE_O0),.C(CLK),.CE(PCI_CE));

IOBUF_PCI33_5 XPCI_PAR      (.O(PAR_I),.IO(PAR),
                             .I(PAR_OUT),.T(OE_PAR_N));
// output flipflops
FDE XPCI_PAROQ (.Q(PAR_OUT),.D(PAR_O),.C(CLK),.CE(PCI_CE));

IOBUF_PCI33_5 XPCI_FRAME    (.O(FRAME_I),.IO(FRAME_N),
                             .I(FRAME_O),.T(OE_FRAME_N));

IOBUF_PCI33_5 XPCI_TRDY     (.O(TRDY_I),.IO(TRDY_N),
                             .I(TRDY_O),.T(OE_TRDY_N));

IOBUF_PCI33_5 XPCI_IRDY     (.O(IRDY_I),.IO(IRDY_N),
                             .I(IRDY_O),.T(OE_IRDY_N));

IOBUF_PCI33_5 XPCI_STOP     (.O(STOP_I),.IO(STOP_N),
                             .I(STOP_O),.T(OE_STOP_N));

IOBUF_PCI33_5 XPCI_DEVSEL   (.O(DEVSEL_I),.IO(DEVSEL_N),
                             .I(DEVSEL_O),.T(OE_DEVSEL_N));

IOBUF_PCI33_5 XPCI_PERR     (.O(PERR_I),.IO(PERR_N),
                             .I(PERR_O),.T(OE_PERR_N));

IOBUF_PCI33_5 XPCI_SERR     (.O(SERR_I),.IO(SERR_N),
                             .I( 1'b0 ),.T(OE_SERR_N));
// outputs
OBUFT_PCI33_5 XPCI_REQ      (.O(REQ_N),.T(OE_REQ_N),.I(REQ_O));
OBUFT_PCI33_5 XPCI_INTA     (.O(INTA_N),.T(OE_INTA_N),.I( 1'b0 ));
// inputs
IBUF_PCI33_5  XPCI_IDSEL    (.O(IDSEL_I),.I(IDSEL));
IBUF_PCI33_5  XPCI_GNT      (.O(GNT_I),.I(GNT_N));
IBUF_PCI33_5  XPCI_RST      (.O(RST_I),.I(RST_N));

// clock
IBUFG_PCI33_5 XPCI_CKI      (.O(NUB),.I(PCLK));
BUFG XPCI_CKA               (.O(CLK),.I(NUB));
// instantiate our PCI interface implementation
PCI PCI(
	.AD_I({AD31, AD30, AD29, AD28, AD27, AD26, AD25, AD24, AD23, AD22, AD21, AD20, AD19, AD18, AD17, AD16, AD15, AD14, AD13, AD12, AD11, AD10, AD9, AD8, AD7, AD6, AD5, AD4, AD3, AD2, AD1, AD0}),
	.AD_O({AD_O31, AD_O30, AD_O29, AD_O28, AD_O27, AD_O26, AD_O25, AD_O24, AD_O23, AD_O22, AD_O21, AD_O20, AD_O19, AD_O18, AD_O17, AD_O16, AD_O15, AD_O14, AD_O13, AD_O12, AD_O11, AD_O10, AD_O9, AD_O8, AD_O7, AD_O6, AD_O5, AD_O4, AD_O3, AD_O2, AD_O1, AD_O0}),
	.OE_AD_N({OE_AD3_N, OE_AD2_N, OE_AD1_N, OE_AD0_N}),
   .CBE_I({CBE3, CBE2, CBE1, CBE0}),
   .CBE_O({CBE_O3, CBE_O2, CBE_O1, CBE_O0}),
	.OE_CBE_N(OE_CBE_N),
	.PAR_I(PAR_I),
	.PAR_O(PAR_O),
	.OE_PAR_N(OE_PAR_N),
	.FRAME_I(FRAME_I),
	.FRAME_O(FRAME_O),
	.OE_FRAME_N(OE_FRAME_N),
	.TRDY_I(TRDY_I),
	.TRDY_O(TRDY_O),
	.OE_TRDY_N(OE_TRDY_N),
	.IRDY_I(IRDY_I),
	.IRDY_O(IRDY_O),
	.OE_IRDY_N(OE_IRDY_N),
	.STOP_I(STOP_I),
	.STOP_O(STOP_O),
	.OE_STOP_N(OE_STOP_N),
	.DEVSEL_I(DEVSEL_I),
	.DEVSEL_O(DEVSEL_O),
	.OE_DEVSEL_N(OE_DEVSEL_N),
	.IDSEL_I(IDSEL_I),
	.PERR_I(PERR_I),
	.PERR_O(PERR_O),	
	.OE_PERR_N(OE_PERR_N),
	.SERR_I(SERR_I),
	.OE_SERR_N(OE_SERR_N),
	.REQ_O(REQ_O),
	.OE_REQ_N(OE_REQ_N),	
	.GNT_I(GNT_I),
   .CLK(CLK),
	.RST_I(RST_I),
	.RST_O(RST),
	.OE_INTA_N(OE_INTA_N),
   .PING_DONE(PING_DONE),
   .PING_REQ(PING_REQ),
   .PCI_CE(PCI_CE)	
);

endmodule
